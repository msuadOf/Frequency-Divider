module connect (
    input wire i_rst_n,
    output wire o_rst_n
);
assign o_rst_n=i_rst_n;
endmodule //connect